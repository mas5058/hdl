 -----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--Michael Sarlo
--lab 1
--9/1/17
--or gate
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;      

entity or3 is 
  port (
    a       : in std_logic;
    b       : in std_logic;
    c       : in std_logic;
	z       : out std_logic
  );
end or3;

architecture arch of or3 is
begin 
  z  <= (a or b or c);
end arch; 