 -----------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
--Michael Sarlo
--lab 1
--9/1/17
--and gate
---------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;      

entity and2 is 
  port (
    a       : in std_logic;
    b       : in std_logic;
	z       : out std_logic
  );
end and2;

architecture arch of and2 is
begin 
  z  <= (a and b);
end arch; 