blink_rom_inst : blink_rom PORT MAP (
        address     => address_sig,
        clock     => clock_sig,
        q     => q_sig
    );
